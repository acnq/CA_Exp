`include "define.vh"


/**
 * Controller for MIPS 5-stage pipelined CPU.
 * Author: Zhao, Hongyu  <power_zhy@foxmail.com>
 */
module controller (/*AUTOARG*/
	input wire clk,  // main clock
	input wire rst,  // synchronous reset
	// debug
	`ifdef DEBUG
	input wire debug_en,  // debug enable
	input wire debug_step,  // debug step clock
	`endif
	// instruction decode
	input wire [31:0] inst,  // instruction
	output reg [2:0] pc_src,  // how would PC change to next
	output reg imm_ext,  // whether using sign extended to immediate data
	output reg [1:0] exe_a_src,  // data source of operand A for ALU
	output reg [1:0] exe_b_src,  // data source of operand B for ALU
	output reg [3:0] exe_alu_oper,  // ALU operation type
	output reg mem_ren,  // memory read enable signal
	output reg mem_wen,  // memory write enable signal
	output reg [1:0] wb_addr_src,  // address source to write data back to registers
	output reg wb_data_src,  // data source of data being written back to registers
	output reg wb_wen,  // register write enable signal
	output reg unrecognized,  // whether current instruction can not be recognized
	// debug control
	output reg cpu_rst,  // cpu reset signal
	output reg cpu_en  // cpu enable signal
	);
	
	`include "mips_define.vh"
	
	// instruction decode
	always @(*) begin
		pc_src = PC_NEXT;
		imm_ext = 0;
		exe_a_src = EXE_A_RS;
		exe_b_src = EXE_B_RT;
		exe_alu_oper = EXE_ALU_ADD;
		mem_ren = 0;
		mem_wen = 0;
		wb_addr_src = WB_ADDR_RD;
		wb_data_src = WB_DATA_ALU;
		wb_wen = 0;
		unrecognized = 0;
		case (inst[31:26])
			INST_R: begin
				case (inst[5:0])
					R_FUNC_JR: begin
						pc_src = PC_JR;
					end
					R_FUNC_ADD: begin
						exe_alu_oper = EXE_ALU_ADD;
						wb_addr_src = WB_ADDR_RD;
						wb_data_src = WB_DATA_ALU;
						wb_wen = 1;
					end
					R_FUNC_SUB: begin
						exe_alu_oper = EXE_ALU_SUB;//
						wb_addr_src = WB_ADDR_RD;//
						wb_data_src = WB_DATA_ALU;//
						wb_wen = 1;
					end
					R_FUNC_AND: begin
						exe_alu_oper = EXE_ALU_AND;
						wb_addr_src = WB_ADDR_RD;
						wb_data_src = WB_DATA_ALU;
						wb_wen = 1;
					end
					R_FUNC_OR: begin
						exe_alu_oper = EXE_ALU_OR;
						wb_addr_src = WB_ADDR_RD;
						wb_data_src = WB_DATA_ALU;
						wb_wen = 1;
					end
					R_FUNC_SLT: begin
						exe_alu_oper = EXE_ALU_SLT;
						wb_addr_src = WB_ADDR_RD;
						wb_data_src = WB_DATA_ALU;
						wb_wen = 1;
					end
					default: begin
						unrecognized = 1;
					end
				endcase
			end
			INST_J: begin
				pc_src = PC_JUMP;//
			end
			INST_JAL: begin
				pc_src = PC_JUMP;//
				exe_a_src = EXE_A_LINK;//
				exe_b_src = EXE_B_LINK;//
				exe_alu_oper = EXE_ALU_ADD;//
				wb_addr_src = WB_ADDR_LINK;//
				wb_data_src = WB_DATA_ALU;//
				wb_wen = 1;
			end
			INST_BEQ: begin
				pc_src = PC_BEQ;//
				exe_a_src = EXE_A_BRANCH;//
				exe_b_src = EXE_B_BRANCH;//
				exe_alu_oper = EXE_ALU_ADD;//
				imm_ext = 1;
			end
			INST_BNE: begin//add myself
				pc_src = PC_BNE;//
				exe_a_src = EXE_A_BRANCH;//
				exe_b_src = EXE_B_BRANCH;//
				exe_alu_oper = EXE_ALU_ADD;//
				imm_ext = 1;
			end
			INST_ADDI: begin
				imm_ext = 1;
				exe_b_src = EXE_B_IMM;
				exe_alu_oper = EXE_ALU_ADD;
				wb_addr_src = WB_ADDR_RT;
				wb_data_src = WB_DATA_ALU;
				wb_wen = 1;
			end
			INST_ANDI: begin
				imm_ext = 0;//Ϊɶ��0?
				exe_b_src = EXE_B_IMM;//
				exe_alu_oper = EXE_ALU_AND;//
				wb_addr_src = WB_ADDR_RT;//
				wb_data_src = WB_DATA_ALU;//
				wb_wen = 1;//
			end
			INST_ORI: begin
				imm_ext = 0;//Ϊɶ��0?
				exe_b_src = EXE_B_IMM;
				exe_alu_oper = EXE_ALU_OR;
				wb_addr_src = WB_ADDR_RT;
				wb_data_src = WB_DATA_ALU;
				wb_wen = 1;
			end
			INST_LW: begin
				imm_ext = 1;//
				exe_b_src = EXE_B_IMM;//
				exe_alu_oper = EXE_ALU_ADD;//
				mem_ren = 1;//
				wb_addr_src = WB_ADDR_RT;//
				wb_data_src = WB_DATA_MEM;//
				wb_wen = 1;
			end
			INST_SW: begin
				imm_ext = 1;//
				exe_b_src = EXE_B_IMM;//
				exe_alu_oper = EXE_ALU_ADD;//
				mem_wen = 1;//
			end
			default: begin
				unrecognized = 1;
			end
		endcase
	end
	
	// debug control
	`ifdef DEBUG
	reg debug_step_prev;
	
	always @(posedge clk) begin
		debug_step_prev <= debug_step;
	end
	`endif
	
	always @(*) begin
		cpu_rst = 0;
		cpu_en = 1;
		if (rst) begin
			cpu_rst = 1;
		end
		`ifdef DEBUG
		// suspend and step execution
		else if ((debug_en) && ~(~debug_step_prev && debug_step)) begin
			cpu_en = 0;
		end
		`endif
	end
	
endmodule
